//Instruction Register
module IR();
endmodule